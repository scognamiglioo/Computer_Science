/*
Guia_0203
*/
module Guia_0203;
// define data
real x = 0.0;
// decimal
reg [7:0] b = 8'b0000_0000 ; // binary 

// actions
initial
begin : main
$display ( "Guia_0203 - Tests" );

//--------------------------------------------------------------//

b = 8'b00_01_11_01;
$display ( " a = %d,%d%d%d" , b[7:6],b[5:4], b[3:2], b[1:0] );
$display ( "---------------------------------------------- ");


//--------------------------------------------------------------//


x = 0.0;
b = 8'b1001_0100;
$display ( " b = %d,%o%o" , x, b[7:5],b[4:2] );
$display ( "---------------------------------------------- ");

//--------------------------------------------------------------//


b = 8'b00_100110;
$display ( " c = %x,%x", b[7:6],b[5:0] );
$display ( "---------------------------------------------- ");

//--------------------------------------------------------------//


x = 1.0;
b = 8'b1100_1100;
$display ( " d = %d,%o%o" , x, b[7:5],b[4:2] );
$display ( "---------------------------------------------- ");

//--------------------------------------------------------------//


b = 8'b1101_1101;
$display ( " e = %x,%x", b[7:4],b[3:0] );
$display ( "---------------------------------------------- ");

end // main
endmodule // Guia_0203